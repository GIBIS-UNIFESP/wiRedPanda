// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 30 LUTs, 38 FFs, 11 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: display_3bits_counter
// Generated: Fri Sep 26 03:03:40 2025
// Target FPGA: Generic-Small
// Resource Usage: 30/1000 LUTs, 38/1000 FFs, 11/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module display_3bits_counter (
    // ========= Input Ports =========
// DEBUG: Input port: Clock -> input_clock1_1 (Element: Clock)
// DEBUG: Input port: Push Button -> input_push_button2_btn_2 (Element: Push Button)
    input wire input_clock1_1,
    input wire input_push_button2_btn_2,

    // ========= Output Ports =========
// DEBUG: Output port: 7-Segment Display[0] -> output_7_segment_display1_g_middle_3 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[1] -> output_7_segment_display1_f_upper_left_4 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[2] -> output_7_segment_display1_e_lower_left_5 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[3] -> output_7_segment_display1_d_bottom_6 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[4] -> output_7_segment_display1_a_top_7 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[5] -> output_7_segment_display1_b_upper_right_8 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[6] -> output_7_segment_display1_dp_dot_9 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[7] -> output_7_segment_display1_c_lower_right_10 (Element: 7-Segment Display)
    output wire output_7_segment_display1_g_middle_3,
    output wire output_7_segment_display1_f_upper_left_4,
    output wire output_7_segment_display1_e_lower_left_5,
    output wire output_7_segment_display1_d_bottom_6,
    output wire output_7_segment_display1_a_top_7,
    output wire output_7_segment_display1_b_upper_right_8,
    output wire output_7_segment_display1_dp_dot_9,
    output wire output_7_segment_display1_c_lower_right_10
);

    // ========= Internal Signals =========
    wire node_11_0;
    reg t_flip_flop_12_0_0 = 1'b0;
    reg t_flip_flop_13_1_1 = 1'b0;
    wire node_14_0;
    reg t_flip_flop_15_0_0 = 1'b0;
    reg t_flip_flop_16_1_1 = 1'b0;
    wire node_17_0;
    reg t_flip_flop_18_0_0 = 1'b0;
    reg t_flip_flop_19_1_1 = 1'b0;
    wire node_20_0;
    wire node_21_0;
    wire node_22_0;
    wire node_23_0;
    wire node_24_0;
    wire node_25_0;
    wire ic_display_3bits_ic_node_26_0;
    wire ic_display_3bits_ic_or_27_0;
    wire ic_display_3bits_ic_or_28_0;
    wire ic_display_3bits_ic_and_29_0;
    wire ic_display_3bits_ic_or_30_0;
    wire ic_display_3bits_ic_not_31_0;
    wire ic_display_3bits_ic_and_32_0;
    wire ic_display_3bits_ic_and_33_0;
    wire ic_display_3bits_ic_and_34_0;
    wire ic_display_3bits_ic_xnor_35_0;
    wire ic_display_3bits_ic_and_36_0;
    wire ic_display_3bits_ic_or_37_0;
    wire ic_display_3bits_ic_nand_38_0;
    wire ic_display_3bits_ic_or_39_0;
    wire ic_display_3bits_ic_or_40_0;
    wire ic_display_3bits_ic_node_41_0;
    wire ic_display_3bits_ic_node_42_0;
    wire ic_display_3bits_ic_node_43_0;
    wire ic_display_3bits_ic_node_44_0;
    wire ic_display_3bits_ic_node_45_0;
    wire ic_display_3bits_ic_node_46_0;
    wire ic_display_3bits_ic_node_47_0;
    wire ic_display_3bits_ic_node_48_0;
    wire ic_display_3bits_ic_not_49_0;
    wire ic_display_3bits_ic_and_50_0;
    wire ic_display_3bits_ic_and_51_0;
    wire ic_display_3bits_ic_and_52_0;
    wire ic_display_3bits_ic_and_53_0;
    wire ic_display_3bits_ic_node_54_0;
    wire ic_display_3bits_ic_or_55_0;
    wire ic_display_3bits_ic_node_56_0;
    wire ic_display_3bits_ic_node_57_0;
    wire ic_display_3bits_ic_xnor_58_0;
    wire ic_display_3bits_ic_gnd_59_0;
    wire ic_display_3bits_ic_or_60_0;
    wire ic_display_3bits_ic_and_61_0;
    wire ic_display_3bits_ic_not_62_0;
    wire ic_display_3bits_ic_or_63_0;
    wire ic_display_3bits_ic_gnd_64_0;

    // ========= Logic Assignments =========
// DEBUG: Processing 16 top-level elements with topological sorting
// DEBUG: Processing 39 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_59_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_59_0 (Element: GND)
    assign ic_display_3bits_ic_node_26_0 = ic_display_3bits_ic_gnd_59_0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_27_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_28_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_29_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_30_0 = (((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_31_0 = ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_32_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_33_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_34_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_xnor_35_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Xnor
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_36_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_37_0 = ((~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_nand_38_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_39_0 = (((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (1'b0 & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_40_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) | (ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_41_0 = (((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (1'b0 & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_42_0 = ((~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_43_0 = (((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_44_0 = ((~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_45_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) | (ic_display_3bits_ic_gnd_64_0 | 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_46_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) | (ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_59_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_59_0 (Element: GND)
    assign ic_display_3bits_ic_node_47_0 = ic_display_3bits_ic_gnd_59_0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_48_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_49_0 = ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_50_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_51_0 = (1'b0 & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_52_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_53_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_54_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_55_0 = ((~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_64_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_56_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_57_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_xnor_58_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Xnor
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_60_0 = ((ic_display_3bits_ic_gnd_64_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_64_0 | 1'b0) | (ic_display_3bits_ic_gnd_64_0 | 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_61_0 = (~(ic_display_3bits_ic_gnd_64_0 | 1'b0) & (ic_display_3bits_ic_gnd_64_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_62_0 = ~(ic_display_3bits_ic_gnd_64_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_64_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_64_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_63_0 = (ic_display_3bits_ic_gnd_64_0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock1_1' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock1_1 (Element: Clock)
    assign node_25_0 = input_clock1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_16_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_16_1_1 (Element: T-Flip-Flop)
    assign node_24_0 = t_flip_flop_16_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_13_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_13_1_1 (Element: T-Flip-Flop)
    assign node_23_0 = t_flip_flop_13_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock1_1' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock1_1 (Element: Clock)
    assign node_22_0 = input_clock1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_19_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_19_1_1 (Element: T-Flip-Flop)
    assign node_21_0 = t_flip_flop_19_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_19_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_19_1_1 (Element: T-Flip-Flop)
    assign node_20_0 = t_flip_flop_19_1_1; // Node
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button2_btn_2' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button2_btn_2 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_16_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_16_1_1 (Element: T-Flip-Flop)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
    // T FlipFlop: T-Flip-Flop
    always @(posedge t_flip_flop_16_1_1) begin
        begin
            if (input_push_button2_btn_2) begin // toggle
                t_flip_flop_18_0_0 <= t_flip_flop_19_1_1;
                t_flip_flop_19_1_1 <= t_flip_flop_18_0_0;
            end
            // else hold
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button2_btn_2' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button2_btn_2 (Element: Push Button)
    assign node_17_0 = input_push_button2_btn_2; // Node
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button2_btn_2' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button2_btn_2 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: T-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 't_flip_flop_13_1_1' (Element: T-Flip-Flop)
// DEBUG: otherPortName: Final result: t_flip_flop_13_1_1 (Element: T-Flip-Flop)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
    // T FlipFlop: T-Flip-Flop
    always @(posedge t_flip_flop_13_1_1) begin
        begin
            if (input_push_button2_btn_2) begin // toggle
                t_flip_flop_15_0_0 <= t_flip_flop_16_1_1;
                t_flip_flop_16_1_1 <= t_flip_flop_15_0_0;
            end
            // else hold
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button2_btn_2' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button2_btn_2 (Element: Push Button)
    assign node_14_0 = input_push_button2_btn_2; // Node
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button2_btn_2' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button2_btn_2 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock1_1' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock1_1 (Element: Clock)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
// DEBUG: otherPortName: Processing port from element T-Flip-Flop (type 20) (Element: T-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: T-Flip-Flop)
    // T FlipFlop: T-Flip-Flop
    always @(posedge input_clock1_1) begin
        begin
            if (input_push_button2_btn_2) begin // toggle
                t_flip_flop_12_0_0 <= t_flip_flop_13_1_1;
                t_flip_flop_13_1_1 <= t_flip_flop_12_0_0;
            end
            // else hold
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock1_1' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock1_1 (Element: Clock)
    assign node_11_0 = input_clock1_1; // Node

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_g_middle_3 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_f_upper_left_4 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_e_lower_left_5 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_d_bottom_6 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_a_top_7 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_b_upper_right_8 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock1_1' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock1_1 (Element: Clock)
    assign output_7_segment_display1_dp_dot_9 = input_clock1_1; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_c_lower_right_10 = 1'b0; // 7-Segment Display

endmodule // display_3bits_counter

// ====================================================================
// Module display_3bits_counter generation completed successfully
// Elements processed: 16
// Inputs: 2, Outputs: 8
// ====================================================================
