// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: dflipflop2_debug
// Generated: Sun Sep 28 00:41:24 2025
// Target FPGA: Generic-Small
// Resource Usage: 28/1000 LUTs, 36/1000 FFs, 4/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

`timescale 1ns/1ps

module dflipflop2_debug (
    // ========= Input Ports =========
    input wire input_clock1_1,
    input wire input_input_switch2_2,

    // ========= Output Ports =========
    output wire output_led1_0_3,
    output wire output_led2_0_4
);

    // ========= Logic Assignments =========

    // ========= Internal Sequential Register =========
    reg output_led1_0_3_behavioral_reg = 1'b0; // Internal sequential register

    // ========= Behavioral Sequential Logic (replaces gate-level feedback) =========
    // Industry-standard behavioral sequential logic
    always @(posedge input_clock1_1) begin
begin // Synchronous operation
            output_led1_0_3_behavioral_reg <= input_input_switch2_2;
        end
    end


    // ========= Output Assignments =========
    // ========= Internal Signals =========

    // ========= Logic Assignments =========
    assign output_led1_0_3 = output_led1_0_3_behavioral_reg; // Connect behavioral register to output
    assign output_led2_0_4 = ~output_led1_0_3_behavioral_reg; // Complementary output
    assign output_led1_0_3 = seq_d_flip_flop_5_0_q; // LED
    assign output_led2_0_4 = ~((input_input_switch2_2 & ~input_clock1_1 & ~(1'b0 & input_clock1_1 & input_input_switch2_2)) & input_clock1_1 & ~(1'b0 & ~(input_clock1_1 & (input_input_switch2_2 & ~input_clock1_1 & 1'b0) & input_clock1_1 & input_input_switch2_2))); // LED


    // ========= ULTRATHINK FINAL SCAN: Diagnostic Information =========
    // ULTRATHINK DEBUG: Found 0 potentially undeclared variables
    // ULTRATHINK DEBUG: Already declared variables count: 2
    // ULTRATHINK DEBUG: Scanned content size: 518 characters
    // ULTRATHINK DEBUG: No additional variables found to declare

endmodule // dflipflop2_debug

// ====================================================================
// Module dflipflop2_debug generation completed successfully
// Elements processed: 24
// Inputs: 2, Outputs: 2
// ====================================================================
