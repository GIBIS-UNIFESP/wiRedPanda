// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 45 LUTs, 74 FFs, 8 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: sequential_debug
// Generated: Fri Sep 26 03:08:01 2025
// Target FPGA: Generic-Small
// Resource Usage: 45/1000 LUTs, 74/1000 FFs, 8/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module sequential_debug (
    // ========= Input Ports =========
// DEBUG: Input port: Push Button -> input_push_button1_reset_1 (Element: Push Button)
// DEBUG: Input port: Clock -> input_clock2_slow_clk_2 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock3_fast_clk_3 (Element: Clock)
    input wire input_push_button1_reset_1,
    input wire input_clock2_slow_clk_2,
    input wire input_clock3_fast_clk_3,

    // ========= Output Ports =========
// DEBUG: Output port: LED[0] -> output_led1_load_shift_0_4 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led2_l1_0_5 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led3_l3_0_6 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led4_l2_0_7 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led5_l0_0_8 (Element: LED)
    output wire output_led1_load_shift_0_4,
    output wire output_led2_l1_0_5,
    output wire output_led3_l3_0_6,
    output wire output_led4_l2_0_7,
    output wire output_led5_l0_0_8
);

    // ========= Internal Signals =========
    wire not_9_0;
    wire node_10_0;
    wire node_11_0;
    reg jk_flip_flop_12_0_0 = 1'b0;
    reg jk_flip_flop_13_1_1 = 1'b0;
    wire node_14_0;
    reg jk_flip_flop_15_0_0 = 1'b0;
    reg jk_flip_flop_16_1_1 = 1'b0;
    wire node_17_0;
    reg jk_flip_flop_18_0_0 = 1'b0;
    reg jk_flip_flop_19_1_1 = 1'b0;
    wire node_20_0;
    reg jk_flip_flop_21_0_0 = 1'b0;
    reg jk_flip_flop_22_1_1 = 1'b0;
    wire node_23_0;
    wire node_24_0;
    wire node_25_0;
    wire node_26_0;
    wire node_27_0;
    wire node_28_0;
    wire node_29_0;
    wire ic_serialize_ic_node_30_0;
    wire ic_serialize_ic_node_31_0;
    wire ic_serialize_ic_node_32_0;
    wire ic_serialize_ic_node_33_0;
    wire ic_serialize_ic_node_34_0;
    wire ic_serialize_ic_node_35_0;
    wire ic_serialize_ic_node_36_0;
    wire ic_serialize_ic_node_37_0;
    wire ic_serialize_ic_node_38_0;
    wire ic_serialize_ic_node_39_0;
    wire ic_serialize_ic_node_40_0;
    wire ic_serialize_ic_node_41_0;
    wire ic_serialize_ic_node_42_0;
    wire ic_serialize_ic_node_43_0;
    wire ic_serialize_ic_node_44_0;
    wire ic_serialize_ic_node_45_0;
    wire ic_serialize_ic_node_46_0;
    wire ic_serialize_ic_and_47_0;
    wire ic_serialize_ic_node_48_0;
    wire ic_serialize_ic_not_49_0;
    wire ic_serialize_ic_and_50_0;
    wire ic_serialize_ic_or_51_0;
    wire ic_serialize_ic_and_52_0;
    reg ic_serialize_ic_d_flip_flop_53_0_0 = 1'b0;
    reg ic_serialize_ic_d_flip_flop_54_1_1 = 1'b0;
    wire ic_serialize_ic_and_55_0;
    wire ic_serialize_ic_or_56_0;
    reg ic_serialize_ic_d_flip_flop_57_0_0 = 1'b0;
    reg ic_serialize_ic_d_flip_flop_58_1_1 = 1'b0;
    wire ic_serialize_ic_and_59_0;
    reg ic_serialize_ic_d_flip_flop_60_0_0 = 1'b0;
    reg ic_serialize_ic_d_flip_flop_61_1_1 = 1'b0;
    wire ic_serialize_ic_node_62_0;
    wire ic_serialize_ic_node_63_0;
    wire ic_serialize_ic_node_64_0;
    wire ic_serialize_ic_node_65_0;
    wire ic_serialize_ic_and_66_0;
    reg ic_serialize_ic_d_flip_flop_67_0_0 = 1'b0;
    reg ic_serialize_ic_d_flip_flop_68_1_1 = 1'b0;
    wire ic_serialize_ic_and_69_0;
    wire ic_serialize_ic_or_70_0;
    wire ic_serialize_ic_node_71_0;
    wire node_72_0;
    wire not_73_0;
    wire node_74_0;
    wire node_75_0;
    wire and_76_0;
    wire node_77_0;
    reg ic_register_ic_d_flip_flop_78_0_0 = 1'b0;
    reg ic_register_ic_d_flip_flop_79_1_1 = 1'b0;
    wire ic_register_ic_node_80_0;
    wire ic_register_ic_node_81_0;
    reg ic_register_ic_d_flip_flop_82_0_0 = 1'b0;
    reg ic_register_ic_d_flip_flop_83_1_1 = 1'b0;
    wire ic_register_ic_node_84_0;
    reg ic_register_ic_d_flip_flop_85_0_0 = 1'b0;
    reg ic_register_ic_d_flip_flop_86_1_1 = 1'b0;
    wire ic_register_ic_node_87_0;
    wire ic_register_ic_node_88_0;
    wire ic_register_ic_node_89_0;
    wire ic_register_ic_node_90_0;
    wire ic_register_ic_node_91_0;
    wire ic_register_ic_node_92_0;
    wire ic_register_ic_node_93_0;
    reg ic_register_ic_d_flip_flop_94_0_0 = 1'b0;
    reg ic_register_ic_d_flip_flop_95_1_1 = 1'b0;
    wire node_96_0;
    wire and_97_0;
    wire and_98_0;
    wire and_99_0;
    wire and_100_0;

    // ========= Logic Assignments =========
// DEBUG: Processing 38 top-level elements with topological sorting
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign and_100_0 = (1'b0 & input_clock2_slow_clk_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign and_99_0 = (1'b0 & input_clock2_slow_clk_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign and_98_0 = (1'b0 & input_clock2_slow_clk_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign and_97_0 = (1'b0 & input_clock2_slow_clk_2); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_96_0 = input_clock2_slow_clk_2; // Node
// DEBUG: Processing 14 IC internal elements without topological sorting
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_register_ic_d_flip_flop_78_0_0, secondOut=ic_register_ic_d_flip_flop_79_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_85_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_85_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ic_register_ic_d_flip_flop_85_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_register_ic_d_flip_flop_78_0_0 <= ic_register_ic_d_flip_flop_85_0_0;
            ic_register_ic_d_flip_flop_79_1_1 <= ~ic_register_ic_d_flip_flop_85_0_0;
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_80_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_81_0 = 1'b0; // Node
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_register_ic_d_flip_flop_82_0_0, secondOut=ic_register_ic_d_flip_flop_83_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_78_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_78_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ic_register_ic_d_flip_flop_78_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_register_ic_d_flip_flop_82_0_0 <= ic_register_ic_d_flip_flop_78_0_0;
            ic_register_ic_d_flip_flop_83_1_1 <= ~ic_register_ic_d_flip_flop_78_0_0;
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_94_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_94_0_0 (Element: D-Flip-Flop)
    assign ic_register_ic_node_84_0 = ic_register_ic_d_flip_flop_94_0_0; // Node
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_register_ic_d_flip_flop_85_0_0, secondOut=ic_register_ic_d_flip_flop_86_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_94_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_94_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ic_register_ic_d_flip_flop_94_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_register_ic_d_flip_flop_85_0_0 <= ic_register_ic_d_flip_flop_94_0_0;
            ic_register_ic_d_flip_flop_86_1_1 <= ~ic_register_ic_d_flip_flop_94_0_0;
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_87_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_78_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_78_0_0 (Element: D-Flip-Flop)
    assign ic_register_ic_node_88_0 = ic_register_ic_d_flip_flop_78_0_0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_82_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_82_0_0 (Element: D-Flip-Flop)
    assign ic_register_ic_node_89_0 = ic_register_ic_d_flip_flop_82_0_0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_90_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_register_ic_d_flip_flop_85_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_register_ic_d_flip_flop_85_0_0 (Element: D-Flip-Flop)
    assign ic_register_ic_node_91_0 = ic_register_ic_d_flip_flop_85_0_0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_92_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_register_ic_node_93_0 = 1'b0; // Node
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_register_ic_d_flip_flop_94_0_0, secondOut=ic_register_ic_d_flip_flop_95_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = 1'b0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_register_ic_d_flip_flop_94_0_0 <= 1'b0;
            ic_register_ic_d_flip_flop_95_1_1 <= ~1'b0;
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_77_0 = input_clock2_slow_clk_2; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock3_fast_clk_3' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock3_fast_clk_3 (Element: Clock)
    assign and_76_0 = (~1'b0 & input_clock3_fast_clk_3); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_75_0 = input_clock2_slow_clk_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock3_fast_clk_3' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock3_fast_clk_3 (Element: Clock)
    assign node_74_0 = input_clock3_fast_clk_3; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign not_73_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_72_0 = input_clock2_slow_clk_2; // Node
// DEBUG: Processing 38 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_30_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_31_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_32_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_33_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_34_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_35_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_36_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_37_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_38_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_39_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_40_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_41_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_42_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_43_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_44_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_45_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_46_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_53_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_53_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_and_47_0 = (~1'b1 & ic_serialize_ic_d_flip_flop_53_0_0); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_53_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_53_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_node_48_0 = (~1'b1 & ic_serialize_ic_d_flip_flop_53_0_0); // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_not_49_0 = ~1'b1; // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_57_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_57_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_and_50_0 = (~1'b1 & ic_serialize_ic_d_flip_flop_57_0_0); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_57_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_57_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_or_51_0 = ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_57_0_0)); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_and_52_0 = (1'b1 & 1'b1); // And
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_serialize_ic_d_flip_flop_53_0_0, secondOut=ic_serialize_ic_d_flip_flop_54_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_57_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_57_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_57_0_0)) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_serialize_ic_d_flip_flop_53_0_0 <= ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_57_0_0));
            ic_serialize_ic_d_flip_flop_54_1_1 <= ~((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_57_0_0));
        end
    end

// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_and_55_0 = (1'b1 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_60_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_60_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_or_56_0 = ((1'b1 & 1'b0) | (~1'b1 & ic_serialize_ic_d_flip_flop_60_0_0)); // Or
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_serialize_ic_d_flip_flop_57_0_0, secondOut=ic_serialize_ic_d_flip_flop_58_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_60_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_60_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ((1'b1 & 1'b0) | (~1'b1 & ic_serialize_ic_d_flip_flop_60_0_0)) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_serialize_ic_d_flip_flop_57_0_0 <= ((1'b1 & 1'b0) | (~1'b1 & ic_serialize_ic_d_flip_flop_60_0_0));
            ic_serialize_ic_d_flip_flop_58_1_1 <= ~((1'b1 & 1'b0) | (~1'b1 & ic_serialize_ic_d_flip_flop_60_0_0));
        end
    end

// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_60_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_60_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_and_59_0 = (~1'b1 & ic_serialize_ic_d_flip_flop_60_0_0); // And
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_serialize_ic_d_flip_flop_60_0_0, secondOut=ic_serialize_ic_d_flip_flop_61_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_67_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_67_0_0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_67_0_0)) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_serialize_ic_d_flip_flop_60_0_0 <= ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_67_0_0));
            ic_serialize_ic_d_flip_flop_61_1_1 <= ~((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_67_0_0));
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_62_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_63_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_64_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_65_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_67_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_67_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_and_66_0 = (~1'b1 & ic_serialize_ic_d_flip_flop_67_0_0); // And
// DEBUG: generateSequentialLogic: Processing DFlipFlop D-Flip-Flop (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: firstOut=ic_serialize_ic_d_flip_flop_67_0_0, secondOut=ic_serialize_ic_d_flip_flop_68_1_1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting data signal from input port 0 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: data signal = 1'b0 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clock signal from input port 1 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: DFlipFlop D-Flip-Flop: CLOCK signal = 1'b0 (THIS IS CRITICAL!) (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting preset signal from input port 2 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: preset signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Getting clear signal from input port 3 (Element: D-Flip-Flop)
// DEBUG: otherPortName: Processing port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: clear signal = 1'b1 (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Building sensitivity list with clock=1'b0 (Element: D-Flip-Flop)
// DEBUG: WARNING: DFlipFlop D-Flip-Flop clock is constant 1'b0, this will cause syntax error! (Element: D-Flip-Flop)
// DEBUG: DFlipFlop D-Flip-Flop: Added 'posedge 1'b0' to sensitivity list (Element: D-Flip-Flop)
    // D FlipFlop: D-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            ic_serialize_ic_d_flip_flop_67_0_0 <= 1'b0;
            ic_serialize_ic_d_flip_flop_68_1_1 <= ~1'b0;
        end
    end

// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_and_69_0 = (1'b1 & 1'b1); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element D-Flip-Flop (type 17) (Element: D-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: D-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'ic_serialize_ic_d_flip_flop_67_0_0' (Element: D-Flip-Flop)
// DEBUG: otherPortName: Final result: ic_serialize_ic_d_flip_flop_67_0_0 (Element: D-Flip-Flop)
    assign ic_serialize_ic_or_70_0 = ((1'b1 & 1'b1) | (~1'b1 & ic_serialize_ic_d_flip_flop_67_0_0)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_serialize_ic_node_71_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock3_fast_clk_3' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock3_fast_clk_3 (Element: Clock)
    assign node_29_0 = input_clock3_fast_clk_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_28_0 = input_clock2_slow_clk_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_22_1_1' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_22_1_1 (Element: JK-Flip-Flop)
    assign node_27_0 = jk_flip_flop_22_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_19_1_1' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_19_1_1 (Element: JK-Flip-Flop)
    assign node_26_0 = jk_flip_flop_19_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_16_1_1' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_16_1_1 (Element: JK-Flip-Flop)
    assign node_25_0 = jk_flip_flop_16_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_13_1_1' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_13_1_1 (Element: JK-Flip-Flop)
    assign node_24_0 = jk_flip_flop_13_1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign node_23_0 = input_clock2_slow_clk_2; // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_18_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_18_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_18_0_0 or posedge input_push_button1_reset_1) begin
        if (input_push_button1_reset_1) begin
            jk_flip_flop_21_0_0 <= 1'b1;
            jk_flip_flop_22_1_1 <= 1'b0;
        end else begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_21_0_0 <= 1'b0; jk_flip_flop_22_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_21_0_0 <= 1'b1; jk_flip_flop_22_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_21_0_0 <= jk_flip_flop_22_1_1; jk_flip_flop_22_1_1 <= jk_flip_flop_21_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign node_20_0 = ~input_push_button1_reset_1; // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_15_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_15_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_15_0_0 or posedge input_push_button1_reset_1) begin
        if (input_push_button1_reset_1) begin
            jk_flip_flop_18_0_0 <= 1'b1;
            jk_flip_flop_19_1_1 <= 1'b0;
        end else begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_18_0_0 <= 1'b0; jk_flip_flop_19_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_18_0_0 <= 1'b1; jk_flip_flop_19_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_18_0_0 <= jk_flip_flop_19_1_1; jk_flip_flop_19_1_1 <= jk_flip_flop_18_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign node_17_0 = ~input_push_button1_reset_1; // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_12_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_12_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_12_0_0 or posedge input_push_button1_reset_1) begin
        if (input_push_button1_reset_1) begin
            jk_flip_flop_15_0_0 <= 1'b1;
            jk_flip_flop_16_1_1 <= 1'b0;
        end else begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_15_0_0 <= 1'b0; jk_flip_flop_16_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_15_0_0 <= 1'b1; jk_flip_flop_16_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_15_0_0 <= jk_flip_flop_16_1_1; jk_flip_flop_16_1_1 <= jk_flip_flop_15_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign node_14_0 = ~input_push_button1_reset_1; // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge input_clock2_slow_clk_2 or posedge input_push_button1_reset_1) begin
        if (input_push_button1_reset_1) begin
            jk_flip_flop_12_0_0 <= 1'b1;
            jk_flip_flop_13_1_1 <= 1'b0;
        end else begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_12_0_0 <= 1'b0; jk_flip_flop_13_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_12_0_0 <= 1'b1; jk_flip_flop_13_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_12_0_0 <= jk_flip_flop_13_1_1; jk_flip_flop_13_1_1 <= jk_flip_flop_12_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign node_11_0 = ~input_push_button1_reset_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign node_10_0 = ~input_push_button1_reset_1; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Push Button (type 1) (Element: Push Button)
// DEBUG: otherPortName: Checking varMap for final result (Element: Push Button)
// DEBUG: otherPortName: varMap lookup result: 'input_push_button1_reset_1' (Element: Push Button)
// DEBUG: otherPortName: Final result: input_push_button1_reset_1 (Element: Push Button)
    assign not_9_0 = ~input_push_button1_reset_1; // Not

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign output_led1_load_shift_0_4 = input_clock2_slow_clk_2; // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign output_led2_l1_0_5 = (1'b0 & input_clock2_slow_clk_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign output_led3_l3_0_6 = (1'b0 & input_clock2_slow_clk_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign output_led4_l2_0_7 = (1'b0 & input_clock2_slow_clk_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock2_slow_clk_2' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock2_slow_clk_2 (Element: Clock)
    assign output_led5_l0_0_8 = (1'b0 & input_clock2_slow_clk_2); // LED

endmodule // sequential_debug

// ====================================================================
// Module sequential_debug generation completed successfully
// Elements processed: 38
// Inputs: 3, Outputs: 5
// ====================================================================
