// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 66 LUTs, 0 FFs, 12 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: decoder
// Generated: Fri Sep 26 03:03:38 2025
// Target FPGA: Generic-Small
// Resource Usage: 66/1000 LUTs, 0/1000 FFs, 12/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module decoder (
    // ========= Input Ports =========
// DEBUG: Input port: Input Switch -> input_input_switch1_1 (Element: Input Switch)
// DEBUG: Input port: Input Switch -> input_input_switch2_2 (Element: Input Switch)
// DEBUG: Input port: Input Switch -> input_input_switch3_3 (Element: Input Switch)
    input wire input_input_switch1_1,
    input wire input_input_switch2_2,
    input wire input_input_switch3_3,

    // ========= Output Ports =========
// DEBUG: Output port: LED[0] -> output_led1_0_4 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led2_0_5 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led3_0_6 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led4_0_7 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led5_0_8 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led6_0_9 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led7_0_10 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led8_0_11 (Element: LED)
    output wire output_led1_0_4,
    output wire output_led2_0_5,
    output wire output_led3_0_6,
    output wire output_led4_0_7,
    output wire output_led5_0_8,
    output wire output_led6_0_9,
    output wire output_led7_0_10,
    output wire output_led8_0_11
);

    // ========= Internal Signals =========
    wire node_12_0;
    wire node_13_0;
    wire node_14_0;
    wire not_15_0;
    wire not_16_0;
    wire not_17_0;
    wire node_18_0;
    wire node_19_0;
    wire node_20_0;
    wire node_21_0;
    wire node_22_0;
    wire node_23_0;
    wire node_24_0;
    wire node_25_0;
    wire node_26_0;
    wire node_27_0;
    wire node_28_0;
    wire node_29_0;
    wire node_30_0;
    wire node_31_0;
    wire node_32_0;
    wire node_33_0;
    wire node_34_0;
    wire node_35_0;
    wire node_36_0;
    wire node_37_0;
    wire node_38_0;
    wire node_39_0;
    wire node_40_0;
    wire node_41_0;
    wire and_42_0;
    wire and_43_0;
    wire and_44_0;
    wire and_45_0;
    wire and_46_0;
    wire and_47_0;
    wire and_48_0;
    wire and_49_0;
    wire node_50_0;
    wire node_51_0;
    wire node_52_0;
    wire node_53_0;
    wire node_54_0;
    wire node_55_0;

    // ========= Logic Assignments =========
// DEBUG: Processing 55 top-level elements with topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_55_0 = ~input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_54_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_53_0 = ~input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_52_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_51_0 = ~input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_50_0 = input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_49_0 = (input_input_switch3_3 & input_input_switch1_1 & input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_48_0 = (input_input_switch3_3 & input_input_switch1_1 & ~input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_47_0 = (input_input_switch3_3 & ~input_input_switch1_1 & input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_46_0 = (input_input_switch3_3 & ~input_input_switch1_1 & ~input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_45_0 = (~input_input_switch3_3 & input_input_switch1_1 & input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_44_0 = (~input_input_switch3_3 & input_input_switch1_1 & ~input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign and_43_0 = (~input_input_switch3_3 & ~input_input_switch1_1 & input_input_switch2_2); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign and_42_0 = (~input_input_switch2_2 & ~input_input_switch1_1 & ~input_input_switch3_3); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_41_0 = input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_40_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_39_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_38_0 = ~input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_37_0 = ~input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_36_0 = ~input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_35_0 = input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_34_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_33_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_32_0 = ~input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_31_0 = ~input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_30_0 = ~input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_29_0 = input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_28_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_27_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_26_0 = ~input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_25_0 = ~input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_24_0 = ~input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_23_0 = input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_22_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_21_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_20_0 = ~input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_19_0 = ~input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_18_0 = ~input_input_switch3_3; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign not_17_0 = ~input_input_switch2_2; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign not_16_0 = ~input_input_switch1_1; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign not_15_0 = ~input_input_switch3_3; // Not
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign node_14_0 = input_input_switch2_2; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
    assign node_13_0 = input_input_switch1_1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign node_12_0 = input_input_switch3_3; // Node

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led1_0_4 = (input_input_switch3_3 & input_input_switch1_1 & input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led2_0_5 = (input_input_switch3_3 & input_input_switch1_1 & ~input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led3_0_6 = (input_input_switch3_3 & ~input_input_switch1_1 & input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led4_0_7 = (input_input_switch3_3 & ~input_input_switch1_1 & ~input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led5_0_8 = (~input_input_switch3_3 & input_input_switch1_1 & input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led6_0_9 = (~input_input_switch3_3 & input_input_switch1_1 & ~input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
    assign output_led7_0_10 = (~input_input_switch3_3 & ~input_input_switch1_1 & input_input_switch2_2); // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_3 (Element: Input Switch)
    assign output_led8_0_11 = (~input_input_switch2_2 & ~input_input_switch1_1 & ~input_input_switch3_3); // LED

endmodule // decoder

// ====================================================================
// Module decoder generation completed successfully
// Elements processed: 55
// Inputs: 3, Outputs: 8
// ====================================================================
