// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 49 LUTs, 0 FFs, 12 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: display_3bits
// Generated: Fri Sep 26 03:03:41 2025
// Target FPGA: Generic-Small
// Resource Usage: 49/1000 LUTs, 0/1000 FFs, 12/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module display_3bits (
    // ========= Input Ports =========
// DEBUG: Input port: Input Switch -> input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: Input port: Input Switch -> input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: Input port: Input Switch -> input_input_switch3_p2_3 (Element: Input Switch)
    input wire input_input_switch1_p3_1,
    input wire input_input_switch2_p1_2,
    input wire input_input_switch3_p2_3,

    // ========= Output Ports =========
// DEBUG: Output port: 7-Segment Display[0] -> output_7_segment_display1_g_middle_4 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[1] -> output_7_segment_display1_f_upper_left_5 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[2] -> output_7_segment_display1_e_lower_left_6 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[3] -> output_7_segment_display1_d_bottom_7 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[4] -> output_7_segment_display1_a_top_8 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[5] -> output_7_segment_display1_b_upper_right_9 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[6] -> output_7_segment_display1_dp_dot_10 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[7] -> output_7_segment_display1_c_lower_right_11 (Element: 7-Segment Display)
    output wire output_7_segment_display1_g_middle_4,
    output wire output_7_segment_display1_f_upper_left_5,
    output wire output_7_segment_display1_e_lower_left_6,
    output wire output_7_segment_display1_d_bottom_7,
    output wire output_7_segment_display1_a_top_8,
    output wire output_7_segment_display1_b_upper_right_9,
    output wire output_7_segment_display1_dp_dot_10,
    output wire output_7_segment_display1_c_lower_right_11
);

    // ========= Internal Signals =========
    wire gnd_12_0;
    wire or_13_0;
    wire or_14_0;
    wire or_15_0;
    wire not_16_0;
    wire not_17_0;
    wire not_18_0;
    wire and_19_0;
    wire and_20_0;
    wire and_21_0;
    wire and_22_0;
    wire xnor_23_0;
    wire and_24_0;
    wire and_25_0;
    wire and_26_0;
    wire and_27_0;
    wire and_28_0;
    wire xnor_29_0;
    wire gnd_30_0;
    wire and_31_0;
    wire node_32_0;
    wire or_33_0;
    wire or_34_0;
    wire nand_35_0;
    wire or_36_0;
    wire or_37_0;
    wire or_38_0;
    wire or_39_0;

    // ========= Logic Assignments =========
// DEBUG: Processing 32 top-level elements with topological sorting
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign or_39_0 = ((gnd_12_0 | input_input_switch2_p1_2) ^ ~(gnd_12_0 | input_input_switch1_p3_1) | (gnd_12_0 | input_input_switch3_p2_3)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_38_0 = ((~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1)) | (~(gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3)) | ((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & (gnd_12_0 | input_input_switch1_p3_1))); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_37_0 = (~(gnd_12_0 | input_input_switch2_p1_2) | (gnd_12_0 | input_input_switch3_p2_3) ^ ~(gnd_12_0 | input_input_switch1_p3_1)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_36_0 = (((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3)) | (~(gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3)) | (input_input_switch3_p2_3 & ~(gnd_12_0 | input_input_switch1_p3_1))); // Or
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign nand_35_0 = (gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1); // Nand
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_34_0 = ((~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1))); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_33_0 = (((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | (~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1))); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_30_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_30_0 (Element: GND)
    assign node_32_0 = gnd_30_0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign and_31_0 = (~(gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3)); // And
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign xnor_29_0 = (gnd_12_0 | input_input_switch2_p1_2) ^ ~(gnd_12_0 | input_input_switch1_p3_1); // Xnor
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_28_0 = (~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_27_0 = (~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_26_0 = (input_input_switch3_p2_3 & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_25_0 = ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & (gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_24_0 = ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign xnor_23_0 = (gnd_12_0 | input_input_switch3_p2_3) ^ ~(gnd_12_0 | input_input_switch1_p3_1); // Xnor
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_22_0 = (~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_21_0 = ((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign and_20_0 = ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign and_19_0 = ((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)); // And
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign not_18_0 = ~(gnd_12_0 | input_input_switch3_p2_3); // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign not_17_0 = ~(gnd_12_0 | input_input_switch1_p3_1); // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
    assign not_16_0 = ~(gnd_12_0 | input_input_switch2_p1_2); // Not
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
    assign or_15_0 = (gnd_12_0 | input_input_switch2_p1_2); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign or_14_0 = (gnd_12_0 | input_input_switch3_p2_3); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign or_13_0 = (gnd_12_0 | input_input_switch1_p3_1); // Or

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_g_middle_4 = (((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3)) | (~(gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3)) | (input_input_switch3_p2_3 & ~(gnd_12_0 | input_input_switch1_p3_1))); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_f_upper_left_5 = ((~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1))); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_e_lower_left_6 = (((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | (~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1))); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_d_bottom_7 = ((~(gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch1_p3_1)) | (~(gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3)) | ((gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1)) | ((gnd_12_0 | input_input_switch2_p1_2) & ~(gnd_12_0 | input_input_switch3_p2_3) & (gnd_12_0 | input_input_switch1_p3_1))); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
    assign output_7_segment_display1_a_top_8 = ((gnd_12_0 | input_input_switch2_p1_2) ^ ~(gnd_12_0 | input_input_switch1_p3_1) | (gnd_12_0 | input_input_switch3_p2_3)); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_b_upper_right_9 = (~(gnd_12_0 | input_input_switch2_p1_2) | (gnd_12_0 | input_input_switch3_p2_3) ^ ~(gnd_12_0 | input_input_switch1_p3_1)); // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_30_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_30_0 (Element: GND)
    assign output_7_segment_display1_dp_dot_10 = gnd_30_0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch2_p1_2' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch2_p1_2 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch3_p2_3' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch3_p2_3 (Element: Input Switch)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'gnd_12_0' (Element: GND)
// DEBUG: otherPortName: Final result: gnd_12_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Input Switch (type 2) (Element: Input Switch)
// DEBUG: otherPortName: Checking varMap for final result (Element: Input Switch)
// DEBUG: otherPortName: varMap lookup result: 'input_input_switch1_p3_1' (Element: Input Switch)
// DEBUG: otherPortName: Final result: input_input_switch1_p3_1 (Element: Input Switch)
    assign output_7_segment_display1_c_lower_right_11 = (gnd_12_0 | input_input_switch2_p1_2) & (gnd_12_0 | input_input_switch3_p2_3) & ~(gnd_12_0 | input_input_switch1_p3_1); // 7-Segment Display

endmodule // display_3bits

// ====================================================================
// Module display_3bits generation completed successfully
// Elements processed: 32
// Inputs: 3, Outputs: 8
// ====================================================================
