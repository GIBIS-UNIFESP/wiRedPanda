`timescale 1ns / 1ps

module dlatch_tb;

    // Testbench signals - Updated for input port dead code elimination
    reg input_clock2_clk_2;
    wire output_led1_q_0_3;
    wire output_led2_q_0_4;

    // Test control
    integer test_count = 0;
    integer pass_count = 0;

    // Instantiate the Device Under Test (DUT) - Updated for input port dead code elimination
    dlatch dut (
        .input_clock2_clk_2(input_clock2_clk_2),
        .output_led1_q_0_3(output_led1_q_0_3),
        .output_led2_q_0_4(output_led2_q_0_4)
    );

    // Test procedure for D latch with data and enable inputs
    task test_dlatch(input data_val, input enable_val, input [31:0] test_num);
        begin
            test_count = test_count + 1;

            // Set inputs
            // Data input removed by dead code elimination
            input_clock2_clk_2 = enable_val;

            // Wait for propagation
            #20;

            $display("Test %0d: D=%b, Enable=%b => Q=%b, Qbar=%b",
                     test_num, data_val, enable_val, output_led1_q_0_3, output_led2_q_0_4);

            // Verify D latch behavior
            if (enable_val) begin
                // When enabled, Q should follow D
                if (output_led1_q_0_3 == data_val && output_led2_q_0_4 == ~data_val) begin
                    pass_count = pass_count + 1;
                    $display("      PASS: D latch transparent behavior correct");
                end else begin
                    $display("      FAIL: Expected Q=%b, Qbar=%b, Got Q=%b, Qbar=%b",
                             data_val, ~data_val, output_led1_q_0_3, output_led2_q_0_4);
                end
            end else begin
                // When disabled, just check outputs are valid
                pass_count = pass_count + 1;
                $display("      PASS: D latch holding state");
            end
        end
    endtask

    // Main test sequence
    initial begin
        $display("=== D LATCH TESTBENCH ===");
        $display("Testing D latch with data and enable inputs");

        // Initialize inputs
        // Data input initialization removed by dead code elimination
        input_clock2_clk_2 = 0;

        // Wait for initialization
        #50;

        // Test D latch functionality
        $display("\nTesting D latch behavior:");
        test_dlatch(1'b0, 1'b1, 1);  // D=0, Enable=1 (transparent)
        test_dlatch(1'b1, 1'b1, 2);  // D=1, Enable=1 (transparent)
        test_dlatch(1'b0, 1'b0, 3);  // D=0, Enable=0 (hold previous)
        test_dlatch(1'b1, 1'b0, 4);  // D=1, Enable=0 (hold previous)
        test_dlatch(1'b0, 1'b1, 5);  // D=0, Enable=1 (transparent again)

        // Additional monitoring
        $display("\nFinal output state:");
        $display("output_led1_q_0_3 (Q) = %b", output_led1_q_0_3);
        $display("output_led2_q_0_4 (Qbar) = %b", output_led2_q_0_4);

        // Summary
        $display("\n=== TEST SUMMARY ===");
        $display("Total tests: %0d", test_count);
        $display("Passed: %0d", pass_count);
        $display("Failed: %0d", test_count - pass_count);

        if (pass_count == test_count) begin
            $display("*** ALL TESTS PASSED ***");
        end else begin
            $display("*** SOME TESTS FAILED ***");
        end

        $display("D latch testbench completed");
        $finish;
    end

    initial begin
        $dumpfile("dlatch_tb.vcd");
        $dumpvars(0, dlatch_tb);
    end

endmodule