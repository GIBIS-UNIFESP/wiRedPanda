// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 16 LUTs, 38 FFs, 9 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: notes
// Generated: Fri Sep 26 03:03:47 2025
// Target FPGA: Generic-Small
// Resource Usage: 16/1000 LUTs, 38/1000 FFs, 9/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module notes (
    // ========= Input Ports =========
// DEBUG: Input port: Clock -> input_clock1_1 (Element: Clock)
    input wire input_clock1_1,

    // ========= Output Ports =========
// DEBUG: Output port: Buzzer[0] -> output_buzzer1_g6_2 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer2_f6_3 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer3_d6_4 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer4_b7_5 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer5_c6_6 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer6_a7_7 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer7_e6_8 (Element: Buzzer)
// DEBUG: Output port: Buzzer[0] -> output_buzzer8_c7_9 (Element: Buzzer)
    output wire output_buzzer1_g6_2,
    output wire output_buzzer2_f6_3,
    output wire output_buzzer3_d6_4,
    output wire output_buzzer4_b7_5,
    output wire output_buzzer5_c6_6,
    output wire output_buzzer6_a7_7,
    output wire output_buzzer7_e6_8,
    output wire output_buzzer8_c7_9
);

    // ========= Internal Signals =========
    wire ic_dflipflop_ic_node_10_0;
    wire ic_dflipflop_ic_node_11_0;
    wire ic_dflipflop_ic_node_12_0;
    wire ic_dflipflop_ic_node_13_0;
    wire ic_dflipflop_ic_nand_14_0;
    wire ic_dflipflop_ic_node_15_0;
    wire ic_dflipflop_ic_nand_16_0;
    wire ic_dflipflop_ic_not_17_0;
    wire ic_dflipflop_ic_nand_18_0;
    wire ic_dflipflop_ic_nand_19_0;
    wire ic_dflipflop_ic_nand_20_0;
    wire ic_dflipflop_ic_nand_21_0;
    wire ic_dflipflop_ic_node_22_0;
    wire ic_dflipflop_ic_not_23_0;
    wire ic_dflipflop_ic_nand_24_0;
    wire ic_dflipflop_ic_nand_25_0;
    wire ic_dflipflop_ic_node_26_0;
    wire ic_dflipflop_ic_node_27_0;
    wire ic_dflipflop_ic_node_28_0;
    wire ic_dflipflop_ic_not_29_0;
    wire ic_dflipflop_ic_node_30_0;
    wire ic_dflipflop_ic_node_31_0;
    wire ic_dflipflop_ic_node_32_0;
    wire ic_dflipflop_ic_node_33_0;
    wire ic_dflipflop_ic_node_34_0;
    wire ic_jkflipflop_ic_node_35_0;
    wire ic_jkflipflop_ic_node_36_0;
    wire ic_jkflipflop_ic_node_37_0;
    wire ic_jkflipflop_ic_node_38_0;
    wire ic_jkflipflop_ic_node_39_0;
    wire ic_jkflipflop_ic_node_40_0;
    wire ic_jkflipflop_ic_node_41_0;
    wire ic_jkflipflop_ic_node_42_0;
    wire ic_jkflipflop_ic_not_43_0;
    wire ic_jkflipflop_ic_and_44_0;
    wire ic_jkflipflop_ic_node_45_0;
    wire ic_jkflipflop_ic_or_46_0;
    wire ic_jkflipflop_ic_node_47_0;
    wire ic_jkflipflop_ic_node_48_0;
    wire ic_jkflipflop_ic_node_49_0;
    wire ic_jkflipflop_ic_node_50_0;
    wire ic_jkflipflop_ic_and_51_0;
    wire ic_jkflipflop_ic_node_52_0;
    wire ic_jkflipflop_ic_node_53_0;
    reg jk_flip_flop_54_0_0 = 1'b0;
    reg jk_flip_flop_55_1_1 = 1'b0;
    reg jk_flip_flop_56_0_0 = 1'b0;
    reg jk_flip_flop_57_1_1 = 1'b0;
    reg jk_flip_flop_58_0_0 = 1'b0;
    reg jk_flip_flop_59_1_1 = 1'b0;
    wire ic_decoder_ic_node_60_0;
    wire ic_decoder_ic_node_61_0;
    wire ic_decoder_ic_node_62_0;
    wire ic_decoder_ic_node_63_0;
    wire ic_decoder_ic_node_64_0;
    wire ic_decoder_ic_node_65_0;
    wire ic_decoder_ic_node_66_0;
    wire ic_decoder_ic_node_67_0;
    wire ic_decoder_ic_not_68_0;
    wire ic_decoder_ic_not_69_0;
    wire ic_decoder_ic_not_70_0;
    wire ic_decoder_ic_node_71_0;
    wire ic_decoder_ic_node_72_0;
    wire ic_decoder_ic_node_73_0;
    wire ic_decoder_ic_node_74_0;
    wire ic_decoder_ic_node_75_0;
    wire ic_decoder_ic_node_76_0;
    wire ic_decoder_ic_node_77_0;
    wire ic_decoder_ic_node_78_0;
    wire ic_decoder_ic_node_79_0;
    wire ic_decoder_ic_node_80_0;
    wire ic_decoder_ic_node_81_0;
    wire ic_decoder_ic_node_82_0;
    wire ic_decoder_ic_and_83_0;
    wire ic_decoder_ic_and_84_0;
    wire ic_decoder_ic_and_85_0;
    wire ic_decoder_ic_and_86_0;
    wire ic_decoder_ic_and_87_0;
    wire ic_decoder_ic_and_88_0;
    wire ic_decoder_ic_and_89_0;
    wire ic_decoder_ic_and_90_0;
    wire ic_decoder_ic_node_91_0;
    wire ic_decoder_ic_node_92_0;
    wire ic_decoder_ic_node_93_0;
    wire ic_decoder_ic_node_94_0;
    wire ic_decoder_ic_node_95_0;
    wire ic_decoder_ic_node_96_0;
    wire ic_decoder_ic_node_97_0;
    wire ic_decoder_ic_node_98_0;
    wire ic_decoder_ic_node_99_0;
    wire ic_decoder_ic_node_100_0;
    wire ic_decoder_ic_node_101_0;
    wire ic_decoder_ic_node_102_0;
    wire ic_decoder_ic_node_103_0;
    wire ic_decoder_ic_node_104_0;
    wire ic_decoder_ic_node_105_0;
    wire ic_decoder_ic_node_106_0;
    wire ic_decoder_ic_node_107_0;
    wire ic_decoder_ic_node_108_0;
    wire ic_decoder_ic_node_109_0;
    wire ic_decoder_ic_node_110_0;
    wire ic_decoder_ic_node_111_0;
    wire ic_decoder_ic_node_112_0;
    wire ic_decoder_ic_node_113_0;
    wire ic_decoder_ic_node_114_0;

    // ========= Logic Assignments =========
// DEBUG: Processing 14 top-level elements with topological sorting
// DEBUG: Processing 55 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_60_0 = (1'b0 & 1'b0 & 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_61_0 = (1'b0 & 1'b0 & ~1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_62_0 = (1'b0 & ~1'b0 & 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_63_0 = (1'b0 & ~1'b0 & ~1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_64_0 = (~1'b0 & 1'b0 & 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_65_0 = (~1'b0 & 1'b0 & ~1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_66_0 = (~1'b0 & ~1'b0 & 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_67_0 = (~1'b0 & ~1'b0 & ~1'b0); // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_not_68_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_not_69_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_not_70_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_71_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_72_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_73_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_74_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_75_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_76_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_77_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_78_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_79_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_80_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_81_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_82_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_83_0 = (~1'b0 & ~1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_84_0 = (~1'b0 & ~1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_85_0 = (~1'b0 & 1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_86_0 = (~1'b0 & 1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_87_0 = (1'b0 & ~1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_88_0 = (1'b0 & ~1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_89_0 = (1'b0 & 1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_and_90_0 = (1'b0 & 1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_91_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_92_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_93_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_94_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_95_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_96_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_97_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_98_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_99_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_100_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_101_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_102_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_103_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_104_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_105_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_106_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_107_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_108_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_109_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_110_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_111_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_112_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_113_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_decoder_ic_node_114_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_56_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_56_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_56_0_0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_58_0_0 <= 1'b0; jk_flip_flop_59_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_58_0_0 <= 1'b1; jk_flip_flop_59_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_58_0_0 <= jk_flip_flop_59_1_1; jk_flip_flop_59_1_1 <= jk_flip_flop_58_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_54_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_54_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_54_0_0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_56_0_0 <= 1'b0; jk_flip_flop_57_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_56_0_0 <= 1'b1; jk_flip_flop_57_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_56_0_0 <= jk_flip_flop_57_1_1; jk_flip_flop_57_1_1 <= jk_flip_flop_56_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_54_0_0 <= 1'b0; jk_flip_flop_55_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_54_0_0 <= 1'b1; jk_flip_flop_55_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_54_0_0 <= jk_flip_flop_55_1_1; jk_flip_flop_55_1_1 <= jk_flip_flop_54_0_0; end // toggle
            endcase
        end
    end

// DEBUG: Processing 20 IC internal elements without topological sorting
// DEBUG: Processing 25 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_10_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_11_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_12_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_13_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_14_0 = ~(1'b0 & ~1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_16_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_16_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_15_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ~(ic_dflipflop_ic_nand_16_0 & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_16_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_16_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_16_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ~(ic_dflipflop_ic_nand_16_0 & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0)); // Nand
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_17_0 = 1'b0; // Not
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_18_0 = (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_19_0 = ~(1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)); // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_20_0 = (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_21_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_21_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_21_0 = (1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ic_dflipflop_ic_nand_21_0) & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_19_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_19_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_21_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_21_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_22_0 = (1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_19_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ic_dflipflop_ic_nand_21_0) & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_23_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_18_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_18_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_24_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_18_0) & 1'b0 & ~1'b0 & 1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_25_0 = 1'b0 & ~1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_26_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_27_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_28_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_29_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_30_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_31_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_32_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_33_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_34_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_35_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_36_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_37_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_38_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_39_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_40_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_41_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_42_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_not_43_0 = ~1'b1; // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_and_44_0 = (1'b1 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_45_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_or_46_0 = ((1'b0 & ~1'b1) | (1'b1 & 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_47_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_48_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_49_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_50_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_and_51_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_52_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_53_0 = 1'b0; // Node

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer1_g6_2 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer2_f6_3 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer3_d6_4 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer4_b7_5 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer5_c6_6 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer6_a7_7 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer7_e6_8 = 1'b0; // Buzzer
// DEBUG: otherPortName: Processing port from element Buzzer (type 26) (Element: Buzzer)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_buzzer8_c7_9 = 1'b0; // Buzzer

endmodule // notes

// ====================================================================
// Module notes generation completed successfully
// Elements processed: 14
// Inputs: 1, Outputs: 8
// ====================================================================
