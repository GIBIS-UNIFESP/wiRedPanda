// DEBUG: Selected FPGA: Generic-Small (Small generic FPGA (educational))
// DEBUG: Estimated resources: 58 LUTs, 215 FFs, 37 IOs
// ====================================================================
// ======= This Verilog code was generated automatically by wiRedPanda =======
// ====================================================================
//
// Module: ic_debug
// Generated: Fri Sep 26 02:46:48 2025
// Target FPGA: Generic-Small
// Resource Usage: 58/1000 LUTs, 215/1000 FFs, 37/50 IOs
//
// wiRedPanda - Digital Logic Circuit Simulator
// https://github.com/gibis-unifesp/wiredpanda
// ====================================================================

module ic_debug (
    // ========= Input Ports =========
// DEBUG: Input port: Clock -> input_clock1_1 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock2_2 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock3_3 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock4_4 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock5_5 (Element: Clock)
// DEBUG: Input port: Clock -> input_clock6_6 (Element: Clock)
    input wire input_clock1_1,
    input wire input_clock2_2,
    input wire input_clock3_3,
    input wire input_clock4_4,
    input wire input_clock5_5,
    input wire input_clock6_6,

    // ========= Output Ports =========
// DEBUG: Output port: 7-Segment Display[0] -> output_7_segment_display1_g_middle_7 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[1] -> output_7_segment_display1_f_upper_left_8 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[2] -> output_7_segment_display1_e_lower_left_9 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[3] -> output_7_segment_display1_d_bottom_10 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[4] -> output_7_segment_display1_a_top_11 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[5] -> output_7_segment_display1_b_upper_right_12 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[6] -> output_7_segment_display1_dp_dot_13 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[7] -> output_7_segment_display1_c_lower_right_14 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[0] -> output_7_segment_display2_g_middle_15 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[1] -> output_7_segment_display2_f_upper_left_16 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[2] -> output_7_segment_display2_e_lower_left_17 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[3] -> output_7_segment_display2_d_bottom_18 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[4] -> output_7_segment_display2_a_top_19 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[5] -> output_7_segment_display2_b_upper_right_20 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[6] -> output_7_segment_display2_dp_dot_21 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[7] -> output_7_segment_display2_c_lower_right_22 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[0] -> output_7_segment_display3_g_middle_23 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[1] -> output_7_segment_display3_f_upper_left_24 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[2] -> output_7_segment_display3_e_lower_left_25 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[3] -> output_7_segment_display3_d_bottom_26 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[4] -> output_7_segment_display3_a_top_27 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[5] -> output_7_segment_display3_b_upper_right_28 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[6] -> output_7_segment_display3_dp_dot_29 (Element: 7-Segment Display)
// DEBUG: Output port: 7-Segment Display[7] -> output_7_segment_display3_c_lower_right_30 (Element: 7-Segment Display)
// DEBUG: Output port: LED[0] -> output_led4_0_31 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led5_0_32 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led6_0_33 (Element: LED)
// DEBUG: Output port: LED[0] -> output_led7_0_34 (Element: LED)
    output wire output_7_segment_display1_g_middle_7,
    output wire output_7_segment_display1_f_upper_left_8,
    output wire output_7_segment_display1_e_lower_left_9,
    output wire output_7_segment_display1_d_bottom_10,
    output wire output_7_segment_display1_a_top_11,
    output wire output_7_segment_display1_b_upper_right_12,
    output wire output_7_segment_display1_dp_dot_13,
    output wire output_7_segment_display1_c_lower_right_14,
    output wire output_7_segment_display2_g_middle_15,
    output wire output_7_segment_display2_f_upper_left_16,
    output wire output_7_segment_display2_e_lower_left_17,
    output wire output_7_segment_display2_d_bottom_18,
    output wire output_7_segment_display2_a_top_19,
    output wire output_7_segment_display2_b_upper_right_20,
    output wire output_7_segment_display2_dp_dot_21,
    output wire output_7_segment_display2_c_lower_right_22,
    output wire output_7_segment_display3_g_middle_23,
    output wire output_7_segment_display3_f_upper_left_24,
    output wire output_7_segment_display3_e_lower_left_25,
    output wire output_7_segment_display3_d_bottom_26,
    output wire output_7_segment_display3_a_top_27,
    output wire output_7_segment_display3_b_upper_right_28,
    output wire output_7_segment_display3_dp_dot_29,
    output wire output_7_segment_display3_c_lower_right_30,
    output wire output_led4_0_31,
    output wire output_led5_0_32,
    output wire output_led6_0_33,
    output wire output_led7_0_34
);

    // ========= Internal Signals =========
    wire ic_dflipflop_ic_node_35_0;
    wire ic_dflipflop_ic_node_36_0;
    wire ic_dflipflop_ic_node_37_0;
    wire ic_dflipflop_ic_node_38_0;
    wire ic_dflipflop_ic_nand_39_0;
    wire ic_dflipflop_ic_node_40_0;
    wire ic_dflipflop_ic_nand_41_0;
    wire ic_dflipflop_ic_not_42_0;
    wire ic_dflipflop_ic_nand_43_0;
    wire ic_dflipflop_ic_nand_44_0;
    wire ic_dflipflop_ic_nand_45_0;
    wire ic_dflipflop_ic_nand_46_0;
    wire ic_dflipflop_ic_node_47_0;
    wire ic_dflipflop_ic_not_48_0;
    wire ic_dflipflop_ic_nand_49_0;
    wire ic_dflipflop_ic_nand_50_0;
    wire ic_dflipflop_ic_node_51_0;
    wire ic_dflipflop_ic_node_52_0;
    wire ic_dflipflop_ic_node_53_0;
    wire ic_dflipflop_ic_not_54_0;
    wire ic_dflipflop_ic_node_55_0;
    wire ic_dflipflop_ic_node_56_0;
    wire ic_dflipflop_ic_node_57_0;
    wire ic_dflipflop_ic_node_58_0;
    wire ic_dflipflop_ic_node_59_0;
    wire ic_jkflipflop_ic_node_60_0;
    wire ic_jkflipflop_ic_node_61_0;
    wire ic_jkflipflop_ic_node_62_0;
    wire ic_jkflipflop_ic_node_63_0;
    wire ic_jkflipflop_ic_node_64_0;
    wire ic_jkflipflop_ic_node_65_0;
    wire ic_jkflipflop_ic_node_66_0;
    wire ic_jkflipflop_ic_node_67_0;
    wire ic_jkflipflop_ic_not_68_0;
    wire ic_jkflipflop_ic_and_69_0;
    wire ic_jkflipflop_ic_node_70_0;
    wire ic_jkflipflop_ic_or_71_0;
    wire ic_jkflipflop_ic_node_72_0;
    wire ic_jkflipflop_ic_node_73_0;
    wire ic_jkflipflop_ic_node_74_0;
    wire ic_jkflipflop_ic_node_75_0;
    wire ic_jkflipflop_ic_and_76_0;
    wire ic_jkflipflop_ic_node_77_0;
    wire ic_jkflipflop_ic_node_78_0;
    reg jk_flip_flop_79_0_0 = 1'b0;
    reg jk_flip_flop_80_1_1 = 1'b0;
    reg jk_flip_flop_81_0_0 = 1'b0;
    reg jk_flip_flop_82_1_1 = 1'b0;
    reg jk_flip_flop_83_0_0 = 1'b0;
    reg jk_flip_flop_84_1_1 = 1'b0;
    wire ic_input_ic_not_85_0;
    wire ic_input_ic_xor_86_0;
    wire ic_input_ic_or_87_0;
    wire ic_input_ic_and_88_0;
    wire ic_input_ic_node_89_0;
    wire ic_input_ic_node_90_0;
    wire ic_input_ic_node_91_0;
    wire ic_input_ic_node_92_0;
    wire ic_input_ic_node_93_0;
    wire ic_input_ic_node_94_0;
    wire ic_display_4bits_ic_node_95_0;
    wire ic_display_4bits_ic_node_96_0;
    wire ic_display_4bits_ic_node_97_0;
    wire ic_display_4bits_ic_node_98_0;
    wire ic_display_4bits_ic_and_99_0;
    wire ic_display_4bits_ic_node_100_0;
    wire ic_display_4bits_ic_node_101_0;
    wire ic_display_4bits_ic_node_102_0;
    wire ic_display_4bits_ic_node_103_0;
    wire ic_display_4bits_ic_node_104_0;
    wire ic_display_4bits_ic_node_105_0;
    wire ic_display_4bits_ic_node_106_0;
    wire ic_display_4bits_ic_node_107_0;
    wire ic_display_4bits_ic_node_108_0;
    wire ic_display_4bits_ic_node_109_0;
    wire ic_display_4bits_ic_node_110_0;
    wire ic_display_4bits_ic_or_111_0;
    wire ic_display_4bits_ic_or_112_0;
    wire ic_display_4bits_ic_node_113_0;
    wire ic_display_4bits_ic_node_114_0;
    wire ic_display_4bits_ic_node_115_0;
    wire ic_display_4bits_ic_node_116_0;
    wire ic_display_4bits_ic_node_117_0;
    wire ic_display_4bits_ic_node_118_0;
    wire ic_display_4bits_ic_node_119_0;
    wire ic_display_4bits_ic_or_120_0;
    wire ic_display_4bits_ic_or_121_0;
    wire ic_display_4bits_ic_or_122_0;
    wire ic_display_4bits_ic_node_123_0;
    wire ic_display_4bits_ic_node_124_0;
    wire ic_display_4bits_ic_node_125_0;
    wire ic_display_4bits_ic_node_126_0;
    wire ic_display_4bits_ic_node_127_0;
    wire ic_display_4bits_ic_node_128_0;
    wire ic_display_4bits_ic_node_129_0;
    wire ic_display_4bits_ic_node_130_0;
    wire ic_display_4bits_ic_node_131_0;
    wire ic_display_4bits_ic_node_132_0;
    wire ic_display_4bits_ic_node_133_0;
    wire ic_display_4bits_ic_or_134_0;
    wire ic_display_4bits_ic_node_135_0;
    wire ic_display_4bits_ic_node_136_0;
    wire ic_display_4bits_ic_node_137_0;
    wire ic_display_4bits_ic_node_138_0;
    wire ic_display_4bits_ic_or_139_0;
    wire ic_display_4bits_ic_and_140_0;
    wire ic_display_4bits_ic_and_141_0;
    wire ic_display_4bits_ic_and_142_0;
    wire ic_display_4bits_ic_and_143_0;
    wire ic_display_4bits_ic_and_144_0;
    wire ic_display_4bits_ic_and_145_0;
    wire ic_display_4bits_ic_node_146_0;
    wire ic_display_4bits_ic_node_147_0;
    wire ic_display_4bits_ic_and_148_0;
    wire ic_display_4bits_ic_node_149_0;
    wire ic_display_4bits_ic_node_150_0;
    wire ic_display_4bits_ic_and_151_0;
    wire ic_display_4bits_ic_node_152_0;
    wire ic_display_4bits_ic_node_153_0;
    wire ic_display_4bits_ic_node_154_0;
    wire ic_display_4bits_ic_node_155_0;
    wire ic_display_4bits_ic_node_156_0;
    wire ic_display_4bits_ic_node_157_0;
    wire ic_display_4bits_ic_node_158_0;
    wire ic_display_4bits_ic_node_159_0;
    wire ic_display_4bits_ic_node_160_0;
    wire ic_display_4bits_ic_node_161_0;
    wire ic_display_4bits_ic_node_162_0;
    wire ic_display_4bits_ic_node_163_0;
    wire ic_display_4bits_ic_node_164_0;
    wire ic_display_4bits_ic_node_165_0;
    wire ic_display_4bits_ic_node_166_0;
    wire ic_display_4bits_ic_node_167_0;
    wire ic_display_4bits_ic_not_168_0;
    wire ic_display_4bits_ic_not_169_0;
    wire ic_display_4bits_ic_not_170_0;
    wire ic_display_4bits_ic_not_171_0;
    wire ic_display_4bits_ic_node_172_0;
    wire ic_display_4bits_ic_node_173_0;
    wire ic_display_4bits_ic_node_174_0;
    wire ic_display_4bits_ic_node_175_0;
    wire ic_display_4bits_ic_and_176_0;
    wire ic_display_4bits_ic_node_177_0;
    wire ic_display_4bits_ic_node_178_0;
    wire ic_display_4bits_ic_node_179_0;
    wire ic_display_4bits_ic_node_180_0;
    wire ic_display_4bits_ic_node_181_0;
    wire ic_display_4bits_ic_node_182_0;
    wire ic_display_4bits_ic_node_183_0;
    wire ic_display_4bits_ic_node_184_0;
    wire ic_display_4bits_ic_node_185_0;
    wire ic_display_4bits_ic_node_186_0;
    wire ic_display_4bits_ic_node_187_0;
    wire ic_display_4bits_ic_or_188_0;
    wire ic_display_4bits_ic_or_189_0;
    wire ic_display_4bits_ic_node_190_0;
    wire ic_display_4bits_ic_node_191_0;
    wire ic_display_4bits_ic_node_192_0;
    wire ic_display_4bits_ic_node_193_0;
    wire ic_display_4bits_ic_node_194_0;
    wire ic_display_4bits_ic_node_195_0;
    wire ic_display_4bits_ic_node_196_0;
    wire ic_display_4bits_ic_or_197_0;
    wire ic_display_4bits_ic_or_198_0;
    wire ic_display_4bits_ic_or_199_0;
    wire ic_display_4bits_ic_node_200_0;
    wire ic_display_4bits_ic_node_201_0;
    wire ic_display_4bits_ic_node_202_0;
    wire ic_display_4bits_ic_node_203_0;
    wire ic_display_4bits_ic_node_204_0;
    wire ic_display_4bits_ic_node_205_0;
    wire ic_display_4bits_ic_node_206_0;
    wire ic_display_4bits_ic_node_207_0;
    wire ic_display_4bits_ic_node_208_0;
    wire ic_display_4bits_ic_node_209_0;
    wire ic_display_4bits_ic_node_210_0;
    wire ic_display_4bits_ic_or_211_0;
    wire ic_display_4bits_ic_node_212_0;
    wire ic_display_4bits_ic_node_213_0;
    wire ic_display_4bits_ic_node_214_0;
    wire ic_display_4bits_ic_node_215_0;
    wire ic_display_4bits_ic_or_216_0;
    wire ic_display_4bits_ic_and_217_0;
    wire ic_display_4bits_ic_and_218_0;
    wire ic_display_4bits_ic_and_219_0;
    wire ic_display_4bits_ic_and_220_0;
    wire ic_display_4bits_ic_and_221_0;
    wire ic_display_4bits_ic_and_222_0;
    wire ic_display_4bits_ic_node_223_0;
    wire ic_display_4bits_ic_node_224_0;
    wire ic_display_4bits_ic_and_225_0;
    wire ic_display_4bits_ic_node_226_0;
    wire ic_display_4bits_ic_node_227_0;
    wire ic_display_4bits_ic_and_228_0;
    wire ic_display_4bits_ic_node_229_0;
    wire ic_display_4bits_ic_node_230_0;
    wire ic_display_4bits_ic_node_231_0;
    wire ic_display_4bits_ic_node_232_0;
    wire ic_display_4bits_ic_node_233_0;
    wire ic_display_4bits_ic_node_234_0;
    wire ic_display_4bits_ic_node_235_0;
    wire ic_display_4bits_ic_node_236_0;
    wire ic_display_4bits_ic_node_237_0;
    wire ic_display_4bits_ic_node_238_0;
    wire ic_display_4bits_ic_node_239_0;
    wire ic_display_4bits_ic_node_240_0;
    wire ic_display_4bits_ic_node_241_0;
    wire ic_display_4bits_ic_node_242_0;
    wire ic_display_4bits_ic_node_243_0;
    wire ic_display_4bits_ic_node_244_0;
    wire ic_display_4bits_ic_not_245_0;
    wire ic_display_4bits_ic_not_246_0;
    wire ic_display_4bits_ic_not_247_0;
    wire ic_display_4bits_ic_not_248_0;
    wire ic_display_3bits_ic_node_249_0;
    wire ic_display_3bits_ic_or_250_0;
    wire ic_display_3bits_ic_or_251_0;
    wire ic_display_3bits_ic_and_252_0;
    wire ic_display_3bits_ic_or_253_0;
    wire ic_display_3bits_ic_not_254_0;
    wire ic_display_3bits_ic_and_255_0;
    wire ic_display_3bits_ic_and_256_0;
    wire ic_display_3bits_ic_and_257_0;
    wire ic_display_3bits_ic_xnor_258_0;
    wire ic_display_3bits_ic_and_259_0;
    wire ic_display_3bits_ic_or_260_0;
    wire ic_display_3bits_ic_nand_261_0;
    wire ic_display_3bits_ic_or_262_0;
    wire ic_display_3bits_ic_or_263_0;
    wire ic_display_3bits_ic_node_264_0;
    wire ic_display_3bits_ic_node_265_0;
    wire ic_display_3bits_ic_node_266_0;
    wire ic_display_3bits_ic_node_267_0;
    wire ic_display_3bits_ic_node_268_0;
    wire ic_display_3bits_ic_node_269_0;
    wire ic_display_3bits_ic_node_270_0;
    wire ic_display_3bits_ic_node_271_0;
    wire ic_display_3bits_ic_not_272_0;
    wire ic_display_3bits_ic_and_273_0;
    wire ic_display_3bits_ic_and_274_0;
    wire ic_display_3bits_ic_and_275_0;
    wire ic_display_3bits_ic_and_276_0;
    wire ic_display_3bits_ic_node_277_0;
    wire ic_display_3bits_ic_or_278_0;
    wire ic_display_3bits_ic_node_279_0;
    wire ic_display_3bits_ic_node_280_0;
    wire ic_display_3bits_ic_xnor_281_0;
    wire ic_display_3bits_ic_gnd_282_0;
    wire ic_display_3bits_ic_or_283_0;
    wire ic_display_3bits_ic_and_284_0;
    wire ic_display_3bits_ic_not_285_0;
    wire ic_display_3bits_ic_or_286_0;
    wire ic_display_3bits_ic_gnd_287_0;
    reg jk_flip_flop_288_0_0 = 1'b0;
    reg jk_flip_flop_289_1_1 = 1'b0;

    // ========= Logic Assignments =========
// DEBUG: Processing 22 top-level elements with topological sorting
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element Clock (type 9) (Element: Clock)
// DEBUG: otherPortName: Checking varMap for final result (Element: Clock)
// DEBUG: otherPortName: varMap lookup result: 'input_clock6_6' (Element: Clock)
// DEBUG: otherPortName: Final result: input_clock6_6 (Element: Clock)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge input_clock6_6) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_288_0_0 <= 1'b0; jk_flip_flop_289_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_288_0_0 <= 1'b1; jk_flip_flop_289_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_288_0_0 <= jk_flip_flop_289_1_1; jk_flip_flop_289_1_1 <= jk_flip_flop_288_0_0; end // toggle
            endcase
        end
    end

// DEBUG: Processing 39 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_282_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_282_0 (Element: GND)
    assign ic_display_3bits_ic_node_249_0 = ic_display_3bits_ic_gnd_282_0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_250_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_251_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_252_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_253_0 = (((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_254_0 = ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_255_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_256_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_257_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_xnor_258_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Xnor
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_259_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_260_0 = ((~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_nand_261_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_262_0 = (((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (1'b0 & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_263_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) | (ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_264_0 = (((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (1'b0 & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_265_0 = ((~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_266_0 = (((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_267_0 = ((~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_268_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) | (ic_display_3bits_ic_gnd_287_0 | 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_269_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) | (ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_282_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_282_0 (Element: GND)
    assign ic_display_3bits_ic_node_270_0 = ic_display_3bits_ic_gnd_282_0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_271_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_272_0 = ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_273_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_274_0 = (1'b0 & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_275_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_276_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_277_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_278_0 = ((~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0)) | ((ic_display_3bits_ic_gnd_287_0 | 1'b0) & ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_279_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_node_280_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_xnor_281_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Xnor
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xnor)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xnor (type 11) (Element: Xnor)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_283_0 = ((ic_display_3bits_ic_gnd_287_0 | 1'b0) ^ ~(ic_display_3bits_ic_gnd_287_0 | 1'b0) | (ic_display_3bits_ic_gnd_287_0 | 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_and_284_0 = (~(ic_display_3bits_ic_gnd_287_0 | 1'b0) & (ic_display_3bits_ic_gnd_287_0 | 1'b0)); // And
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_not_285_0 = ~(ic_display_3bits_ic_gnd_287_0 | 1'b0); // Not
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element GND (type 13) (Element: GND)
// DEBUG: otherPortName: Checking varMap for final result (Element: GND)
// DEBUG: otherPortName: varMap lookup result: 'ic_display_3bits_ic_gnd_287_0' (Element: GND)
// DEBUG: otherPortName: Final result: ic_display_3bits_ic_gnd_287_0 (Element: GND)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_3bits_ic_or_286_0 = (ic_display_3bits_ic_gnd_287_0 | 1'b0); // Or
// DEBUG: Processing 77 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_172_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_173_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_174_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_175_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_176_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_177_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_178_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_179_0 = (1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_180_0 = (1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_181_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_182_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_183_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_184_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_185_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_186_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_187_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_188_0 = ((1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0 | (~1'b0 & 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_189_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_190_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_191_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_192_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_193_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_194_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_195_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_196_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_197_0 = (1'b0 | ~1'b0 | 1'b1); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_198_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_199_0 = (1'b0 | (~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (~1'b0 & 1'b0) | (1'b1 & (1'b0 & ~1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_200_0 = ((1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0 | (~1'b0 & 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_201_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_202_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_203_0 = (1'b0 | (~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (~1'b0 & 1'b0) | (1'b1 & (1'b0 & ~1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_204_0 = ((1'b0 & 1'b1) | 1'b0 | 1'b0 | (~1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_205_0 = ((1'b0 & 1'b1) | ~1'b0 | (~1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_206_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_207_0 = (1'b0 | ~1'b0 | 1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_208_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_209_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_210_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_211_0 = ((1'b0 & 1'b1) | ~1'b0 | (~1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_212_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_213_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_214_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_215_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_216_0 = ((1'b0 & 1'b1) | 1'b0 | 1'b0 | (~1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_217_0 = (1'b1 & (1'b0 & ~1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_218_0 = (1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_219_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_220_0 = (~1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_221_0 = (1'b0 & 1'b1); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_222_0 = (~1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_223_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_224_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_225_0 = (~1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_226_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_227_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_228_0 = (1'b0 & 1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_229_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_230_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_231_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_232_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_233_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_234_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_235_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_236_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_237_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_238_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_239_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_240_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_241_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_242_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_243_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_244_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_245_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_246_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_247_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_248_0 = ~1'b1; // Not
// DEBUG: Processing 77 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_95_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_96_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_97_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_98_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_99_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_100_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_101_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_102_0 = (1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_103_0 = (1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_104_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_105_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_106_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_107_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_108_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_109_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_110_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_111_0 = ((1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0 | (~1'b0 & 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_112_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_113_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_114_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_115_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_116_0 = (~1'b0 & ~1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_117_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_118_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_119_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_120_0 = (1'b0 | ~1'b0 | 1'b1); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_121_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_122_0 = (1'b0 | (~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (~1'b0 & 1'b0) | (1'b1 & (1'b0 & ~1'b0))); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_123_0 = ((1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0 | (~1'b0 & 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_124_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (1'b0 & ~1'b0) | 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_125_0 = ((~1'b0 & ~1'b1) | (1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_126_0 = (1'b0 | (~1'b0 & ~1'b1) | (1'b0 & ~1'b1) | (~1'b0 & 1'b0) | (1'b1 & (1'b0 & ~1'b0))); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_127_0 = ((1'b0 & 1'b1) | 1'b0 | 1'b0 | (~1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_128_0 = ((1'b0 & 1'b1) | ~1'b0 | (~1'b0 & ~1'b1)); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_129_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_130_0 = (1'b0 | ~1'b0 | 1'b1); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_131_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_132_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_133_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_134_0 = ((1'b0 & 1'b1) | ~1'b0 | (~1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_135_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_136_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_137_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_138_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_or_139_0 = ((1'b0 & 1'b1) | 1'b0 | 1'b0 | (~1'b0 & ~1'b1)); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_140_0 = (1'b1 & (1'b0 & ~1'b0)); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_141_0 = (1'b0 & ~1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_142_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_143_0 = (~1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_144_0 = (1'b0 & 1'b1); // And
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_145_0 = (~1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_146_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_147_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_148_0 = (~1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_149_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_150_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_and_151_0 = (1'b0 & 1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_152_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_153_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_154_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_155_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_156_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_157_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_158_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_159_0 = ~1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_160_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_161_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_162_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_163_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_164_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_165_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_166_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_node_167_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_168_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_169_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_170_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_display_4bits_ic_not_171_0 = ~1'b1; // Not
// DEBUG: Processing 10 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_not_85_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Xor (type 10) (Element: Xor)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xor (type 10) (Element: Xor)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_xor_86_0 = (1'b0 ^ 1'b0); // Xor
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_or_87_0 = (1'b0 | 1'b0); // Or
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_and_88_0 = (1'b0 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_89_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_90_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Xor (type 10) (Element: Xor)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Xor)
// DEBUG: otherPortName: Processing port from element Xor (type 10) (Element: Xor)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Xor (type 10) (Element: Xor)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_91_0 = (1'b0 ^ 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_92_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_93_0 = (1'b0 & 1'b0); // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Or)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_input_ic_node_94_0 = (1'b0 | 1'b0); // Node
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_81_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_81_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_81_0_0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_83_0_0 <= 1'b0; jk_flip_flop_84_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_83_0_0 <= 1'b1; jk_flip_flop_84_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_83_0_0 <= jk_flip_flop_84_1_1; jk_flip_flop_84_1_1 <= jk_flip_flop_83_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_79_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_79_0_0 (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge jk_flip_flop_79_0_0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_81_0_0 <= 1'b0; jk_flip_flop_82_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_81_0_0 <= 1'b1; jk_flip_flop_82_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_81_0_0 <= jk_flip_flop_82_1_1; jk_flip_flop_82_1_1 <= jk_flip_flop_81_0_0; end // toggle
            endcase
        end
    end

// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Processing port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: port has no connections, returning default value (Element: JK-Flip-Flop)
    // JK FlipFlop: JK-Flip-Flop
    always @(posedge 1'b0) begin
        begin
            case ({1'b1, 1'b1})
                2'b00: begin /* hold */ end
                2'b01: begin jk_flip_flop_79_0_0 <= 1'b0; jk_flip_flop_80_1_1 <= 1'b1; end
                2'b10: begin jk_flip_flop_79_0_0 <= 1'b1; jk_flip_flop_80_1_1 <= 1'b0; end
                2'b11: begin jk_flip_flop_79_0_0 <= jk_flip_flop_80_1_1; jk_flip_flop_80_1_1 <= jk_flip_flop_79_0_0; end // toggle
            endcase
        end
    end

// DEBUG: Processing 20 IC internal elements without topological sorting
// DEBUG: Processing 25 IC internal elements without topological sorting
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_35_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_36_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_37_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_38_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_39_0 = ~(1'b0 & ~1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_41_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_41_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_40_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ~(ic_dflipflop_ic_nand_41_0 & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0)); // Node
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_41_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_41_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_41_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ~(ic_dflipflop_ic_nand_41_0 & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0)); // Nand
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_42_0 = 1'b0; // Not
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_43_0 = (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_44_0 = ~(1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)); // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_45_0 = (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_46_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_46_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_46_0 = (1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ic_dflipflop_ic_nand_46_0) & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_44_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_44_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_46_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_46_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_47_0 = (1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ~(ic_dflipflop_ic_nand_44_0 & 1'b0 & ~1'b0 & 1'b0)) & 1'b0 & ic_dflipflop_ic_nand_46_0) & ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0) & 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_48_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Circular dependency detected, checking varMap (Element: Nand)
// DEBUG: otherPortName: varMap result for circular dependency: 'ic_dflipflop_ic_nand_43_0' (Element: Nand)
// DEBUG: otherPortName: Returning varMap result for circular dependency: ic_dflipflop_ic_nand_43_0 (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Nand)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_49_0 = ~(1'b0 & (1'b0 & ~(1'b0 & ~1'b0) & ic_dflipflop_ic_nand_43_0) & 1'b0 & ~1'b0 & 1'b0); // Nand
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Nand (type 7) (Element: Nand)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_nand_50_0 = 1'b0 & ~1'b0; // Nand
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_51_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_52_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_53_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_not_54_0 = ~1'b0; // Not
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_55_0 = ~1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_56_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_57_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_58_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_dflipflop_ic_node_59_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_60_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_61_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_62_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_63_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_64_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_65_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_66_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_67_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_not_68_0 = ~1'b1; // Not
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_and_69_0 = (1'b1 & 1'b0); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_70_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element Or (type 6) (Element: Or)
// DEBUG: otherPortName: Found connected port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: And)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_or_71_0 = ((1'b0 & ~1'b1) | (1'b1 & 1'b0)); // Or
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_72_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_73_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_74_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_node_75_0 = 1'b1; // Node
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
// DEBUG: otherPortName: Processing port from element And (type 5) (Element: And)
// DEBUG: otherPortName: Found connected port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Not)
// DEBUG: otherPortName: Processing port from element Not (type 4) (Element: Not)
// DEBUG: otherPortName: Found connected port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Connected to logic gate, generating expression (Element: Node)
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: port has no connections, returning default value (Element: Node)
    assign ic_jkflipflop_ic_and_76_0 = (1'b0 & ~1'b1); // And
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_77_0 = 1'b0; // Node
// DEBUG: otherPortName: Processing port from element Node (type 23) (Element: Node)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign ic_jkflipflop_ic_node_78_0 = 1'b0; // Node

    // ========= Output Assignments =========
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_g_middle_7 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_f_upper_left_8 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_e_lower_left_9 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_d_bottom_10 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_a_top_11 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_b_upper_right_12 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_dp_dot_13 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display1_c_lower_right_14 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_g_middle_15 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_f_upper_left_16 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_e_lower_left_17 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_d_bottom_18 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_a_top_19 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_b_upper_right_20 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_dp_dot_21 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display2_c_lower_right_22 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_g_middle_23 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_f_upper_left_24 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_e_lower_left_25 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_d_bottom_26 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_a_top_27 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_b_upper_right_28 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_dp_dot_29 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element 7-Segment Display (type 14) (Element: 7-Segment Display)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_7_segment_display3_c_lower_right_30 = 1'b0; // 7-Segment Display
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_led4_0_31 = 1'b0; // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_led5_0_32 = 1'b0; // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element IC (type 22) (Element: IC)
// DEBUG: otherPortName: Checking varMap for final result (Element: IC)
// DEBUG: otherPortName: varMap lookup result: '' (Element: IC)
// DEBUG: otherPortName: varMap empty, returning default value (Element: IC)
    assign output_led6_0_33 = 1'b0; // LED
// DEBUG: otherPortName: Processing port from element LED (type 3) (Element: LED)
// DEBUG: otherPortName: Found connected port from element JK-Flip-Flop (type 18) (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Checking varMap for final result (Element: JK-Flip-Flop)
// DEBUG: otherPortName: varMap lookup result: 'jk_flip_flop_288_0_0' (Element: JK-Flip-Flop)
// DEBUG: otherPortName: Final result: jk_flip_flop_288_0_0 (Element: JK-Flip-Flop)
    assign output_led7_0_34 = jk_flip_flop_288_0_0; // LED

endmodule // ic_debug

// ====================================================================
// Module ic_debug generation completed successfully
// Elements processed: 22
// Inputs: 6, Outputs: 28
// ====================================================================
